module MOV(In1, In2);
input [31:0] In1;
output [31:0] In2;
assign In2 = In1;

endmodule